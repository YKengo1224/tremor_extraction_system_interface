kengo@sirotan.9111:1686189116